// Copyright (c) 2022 W-Mai
// 
// This software is released under the MIT License.
// https://opensource.org/licenses/MIT

`include "../core/defines.v"

module xrv32i(
    input clk,
    input rst,

    input [`InstByteBus]    inst_in,        // 指令输入

    output [`MemAddressBus] inst_addr_out,  // 指令地址输出
);



endmodule
