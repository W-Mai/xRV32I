module pc_reg(
	input wire clk
);



endmodule
